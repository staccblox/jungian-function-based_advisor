module
  initial
    $display("ISXP <-> ENXJ, INXP <-> ESXJ, ISXJ <-> ENXP, INXJ <-> ESXP.");
endmodule
