module software_process_aid;
initial begin
   $display ("Use a SDLC (Waterfall/Agile/etc.) as a process for projects for products, & project size (small/medium/large) for timespan.");
   #10 $finish;
end
endmodule
