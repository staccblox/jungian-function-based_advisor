module software_project_management_aid;
initial begin
   $display ("Use a SDLC as a process for projects for products, & project size for timespan.");
   #10 $finish;
end
endmodule
