module software_process_aid;
initial begin
   $display ("Use a SDLC (Waterfall/Agile/etc.) as a process for projects for products, & project size (small/medium/large) for timespan. ");
   $display ("With regards to process elements, six analysis/design layers are architectural (where), data/class (what), interface (how), procedural (when), component (why), and deployment (who); these may correspond to. ");
   $display ("Diagrams by modeling spaces may be recommended: problem (use case & activity) during planning, solution (class & sequence) during analysis & design, and architectural (component & deployment) during implementation/etc. ");
   #10 $finish;
end
endmodule
